--------------------------------------------------------------------------------
-- Company: 
-- Engineer:
--
-- Create Date:   21:38:40 03/14/2021
-- Design Name:   
-- Module Name:   D:/Tugas/VHDLorsomeshitidk/SAP1nome/MARtb.vhd
-- Project Name:  SAP1nome
-- Target Device:  
-- Tool versions:  
-- Description:   
-- 
-- VHDL Test Bench Created by ISE for module: MAR
-- 
-- Dependencies:
-- 
-- Revision:
-- Revision 0.01 - File Created
-- Additional Comments:
--
-- Notes: 
-- This testbench has been automatically generated using types std_logic and
-- std_logic_vector for the ports of the unit under test.  Xilinx recommends
-- that these types always be used for the top-level I/O of a design in order
-- to guarantee that the testbench will bind correctly to the post-implementation 
-- simulation model.
--------------------------------------------------------------------------------
LIBRARY ieee;
USE ieee.std_logic_1164.ALL;
 
-- Uncomment the following library declaration if using
-- arithmetic functions with Signed or Unsigned values
--USE ieee.numeric_std.ALL;
 
ENTITY MARtb IS
END MARtb;
 
ARCHITECTURE behavior OF MARtb IS 
 
    -- Component Declaration for the Unit Under Test (UUT)
 
    COMPONENT MAR
    PORT(
         CLK : IN  std_logic;
         nLm : IN  std_logic;
         inMAR : IN  std_logic_vector(3 downto 0);
         outMAR : OUT  std_logic_vector(3 downto 0)
        );
    END COMPONENT;
    

   --Inputs
   signal CLK : std_logic := '0';
   signal nLm : std_logic := '0';
   signal inMAR : std_logic_vector(3 downto 0) := (others => '0');

 	--Outputs
   signal outMAR : std_logic_vector(3 downto 0);

   -- Clock period definitions
   constant CLK_period : time := 10 ns;
 
BEGIN
 
	-- Instantiate the Unit Under Test (UUT)
   uut: MAR PORT MAP (
          CLK => CLK,
          nLm => nLm,
          inMAR => inMAR,
          outMAR => outMAR
        );

   -- Clock process definitions
   CLK_process :process
   begin
		CLK <= '0';
		wait for CLK_period/2;
		CLK <= '1';
		wait for CLK_period/2;
   end process;
 

  -- Stimulus process
   stim_proc: process
   begin		
     inMAR <= "0111";
	  nLm <= '1';
	  wait for CLK_period/2;
	  nLm <= '0';
	  wait;
   end process;

END;
